use v5.16

print "Hello World\n"; 

my $name = 'Derek'; 

my ($age,$street) = (40,'123 Main St'); 